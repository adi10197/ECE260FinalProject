// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Please do not spread this code without permission 

`timescale 1ns/1ps

module fullchip_tb;

parameter total_cycle = 8;   // how many streamed Q vectors will be processed
parameter bw = 8;            // Q & K vector bit precision
parameter bw_psum = 2*bw+4;  // partial sum bit precision
parameter pr = 16;           // how many products added in each dot product 
parameter col = 16;           // how many dot product units are equipped

integer qk_file ; // file handler
integer qk_scan_file ; // file handler


integer  captured_data;
integer  weight [col*pr-1:0];
`define NULL 0




integer  K[col-1:0][pr-1:0];
integer  Q[total_cycle-1:0][pr-1:0];
integer  result[total_cycle-1:0][col-1:0];
integer  sum[total_cycle-1:0];
integer  fifo_out[total_cycle-1:0];
integer  result_div[total_cycle-1:0][col-1:0]; 
integer  i,j,k,t,p,q,s,u, m;
integer  result_temp;
integer  div_temp = 20'h004dd;

reg reset = 1;
reg clk = 0;
reg [pr*bw-1:0] mem_in_0, mem_in_1; 
reg ofifo_rd = 0;
wire [16:0] inst; 
reg qmem_rd = 0;
reg qmem_wr = 0; 
reg kmem_rd = 0; 
reg kmem_wr = 0;
reg pmem_rd = 0; 
reg pmem_wr = 0; 
reg execute = 0;
reg load = 0;
reg [3:0] qkmem_add = 0;
reg [3:0] pmem_add = 0;
reg acc0, acc1, div0, div1, canRead_0, canRead_1;

wire [bw_psum*col-1:0] sfp_out;

assign inst[16] = ofifo_rd;
assign inst[15:12] = qkmem_add;
assign inst[11:8]  = pmem_add;
assign inst[7] = execute;
assign inst[6] = load;
assign inst[5] = qmem_rd;
assign inst[4] = qmem_wr;
assign inst[3] = kmem_rd;
assign inst[2] = kmem_wr;
assign inst[1] = pmem_rd;
assign inst[0] = pmem_wr;

reg [bw_psum-1:0] temp5b;
reg [bw_psum+3:0] temp_sum;
wire [bw_psum+3:0] sum_out;
reg [bw_psum*col-1:0] temp16b;
wire [2*bw_psum*col-1:0] chip_out;

fullchip #(.bw(bw), .bw_psum(bw_psum), .col(col), .pr(pr)) fullchip_instance (
      .clk0(clk), 
      .clk1(clk), 
      .mem_in_0(mem_in_0), 
      .mem_in_1(mem_in_1), 
      .inst(inst), 
      .div0(div0), 
      .div1(div1), 
      .acc0(acc0), 
      .acc1(acc1), 
      .reset(reset), 
      .canRead_0(canRead_0), 
      .canRead_1(canRead_1),
      .out(chip_out)
);

initial begin 

  $dumpfile("fullchip_tb.vcd");
  $dumpvars(0,fullchip_tb);



///// Q data txt reading /////

$display("##### Q data txt reading #####");


  qk_file = $fopen("qdata.txt", "r");

  //// To get rid of first 3 lines in data file ////
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);


  for (q=0; q<total_cycle; q=q+1) begin
    for (j=0; j<pr; j=j+1) begin
          qk_scan_file = $fscanf(qk_file, "%d\n", captured_data);
          Q[q][j] = captured_data;
          //$display("%d\n", K[q][j]);
    end
  end
/////////////////////////////////


  for (q=0; q<2; q=q+1) begin
    #0.5 clk = 1'b0;   
    #0.5 clk = 1'b1;   
  end


///// K data txt reading /////

$display("##### K data txt reading #####");

  for (q=0; q<10; q=q+1) begin
    #0.5 clk = 1'b0;   
    #0.5 clk = 1'b1;   
  end
  reset = 0;

  qk_file = $fopen("kdata_core0.txt", "r");

  //// To get rid of first 4 lines in data file ////
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);

  for (q=0; q<col/2; q=q+1) begin
    for (j=0; j<pr; j=j+1) begin
          qk_scan_file = $fscanf(qk_file, "%d\n", captured_data);
          K[q][j] = captured_data;
    end
  end

  qk_file = $fopen("kdata_core1.txt", "r");

  //// To get rid of first 4 lines in data file ////
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);
  qk_scan_file = $fscanf(qk_file, "%s\n", captured_data);

  for (q=col/2; q<col; q=q+1) begin
    for (j=0; j<pr; j=j+1) begin
          qk_scan_file = $fscanf(qk_file, "%d\n", captured_data);
          K[q][j] = captured_data;
    end
  end

/////////////// Estimated result printing /////////////////

$display("##### Estimated multiplication result #####");

  for (t=0; t<total_cycle; t=t+1) begin
     for (q=0; q<col; q=q+1) begin
       result[t][q] = 0;
     end
  end

  for (t=0; t<total_cycle; t=t+1) begin
     for (q=0; q<col; q=q+1) begin
         for (k=0; k<pr; k=k+1) begin
            result[t][q] = result[t][q] + Q[t][k] * K[q][k];
         end
     end
  end  
  for (t=0; t<total_cycle; t=t+1) begin
    sum[t]=0;
     for (q=0; q<col; q=q+1) begin
        if (result[t][q] > 0) begin
          sum[t] = sum[t] + result[t][q];
        end
        else begin
          sum[t] = sum[t] - result[t][q];
        end
     end  
  end

  
  for (t=0; t<total_cycle; t=t+1) begin
     for (q=0; q<col; q=q+1) begin

         result_div[t][q] = (result[t][q]<<8)/sum[t][bw_psum +3:7];
         result_temp = (result[t][q]<<8)/div_temp;
        //  $display("output at %d row and %d column is %h", t, q, result_div[t][q]);
         temp5b = result_div[t][q];
         temp16b = {temp16b[139:0], temp5b};
     end
   
    //  $display("prd @cycle%2d: %40h", t, temp16b);
  end

//////////////////////////////////////////////

///// Qmem writing  /////

$display("##### Qmem writing  #####");

  for (q=0; q<total_cycle; q=q+1) begin

    #0.5 clk = 1'b0;  
    qmem_wr = 1;  if (q>0) qkmem_add = qkmem_add + 1; 
    
    mem_in_0[1*bw-1:0*bw] = Q[q][0];
    mem_in_0[2*bw-1:1*bw] = Q[q][1];
    mem_in_0[3*bw-1:2*bw] = Q[q][2];
    mem_in_0[4*bw-1:3*bw] = Q[q][3];
    mem_in_0[5*bw-1:4*bw] = Q[q][4];
    mem_in_0[6*bw-1:5*bw] = Q[q][5];
    mem_in_0[7*bw-1:6*bw] = Q[q][6];
    mem_in_0[8*bw-1:7*bw] = Q[q][7];
    mem_in_0[9*bw-1:8*bw] = Q[q][8];
    mem_in_0[10*bw-1:9*bw] = Q[q][9];
    mem_in_0[11*bw-1:10*bw] = Q[q][10];
    mem_in_0[12*bw-1:11*bw] = Q[q][11];
    mem_in_0[13*bw-1:12*bw] = Q[q][12];
    mem_in_0[14*bw-1:13*bw] = Q[q][13];
    mem_in_0[15*bw-1:14*bw] = Q[q][14];
    mem_in_0[16*bw-1:15*bw] = Q[q][15];

    mem_in_1[1*bw-1:0*bw] = Q[q][0];
    mem_in_1[2*bw-1:1*bw] = Q[q][1];
    mem_in_1[3*bw-1:2*bw] = Q[q][2];
    mem_in_1[4*bw-1:3*bw] = Q[q][3];
    mem_in_1[5*bw-1:4*bw] = Q[q][4];
    mem_in_1[6*bw-1:5*bw] = Q[q][5];
    mem_in_1[7*bw-1:6*bw] = Q[q][6];
    mem_in_1[8*bw-1:7*bw] = Q[q][7];
    mem_in_1[9*bw-1:8*bw] = Q[q][8];
    mem_in_1[10*bw-1:9*bw] = Q[q][9];
    mem_in_1[11*bw-1:10*bw] = Q[q][10];
    mem_in_1[12*bw-1:11*bw] = Q[q][11];
    mem_in_1[13*bw-1:12*bw] = Q[q][12];
    mem_in_1[14*bw-1:13*bw] = Q[q][13];
    mem_in_1[15*bw-1:14*bw] = Q[q][14];
    mem_in_1[16*bw-1:15*bw] = Q[q][15];

    #0.5 clk = 1'b1;  

  end



  #0.5 clk = 1'b0;  
  qmem_wr = 0; 
  qkmem_add = 0;
  #0.5 clk = 1'b1;  
///////////////////////////////////////////





///// Kmem writing  /////

$display("##### Kmem writing #####");

  for (q=0; q<col/2; q=q+1) begin

    #0.5 clk = 1'b0;  
    kmem_wr = 1; if (q>0) qkmem_add = qkmem_add + 1; 
    
    mem_in_0[1*bw-1:0*bw] = K[q][0];
    mem_in_0[2*bw-1:1*bw] = K[q][1];
    mem_in_0[3*bw-1:2*bw] = K[q][2];
    mem_in_0[4*bw-1:3*bw] = K[q][3];
    mem_in_0[5*bw-1:4*bw] = K[q][4];
    mem_in_0[6*bw-1:5*bw] = K[q][5];
    mem_in_0[7*bw-1:6*bw] = K[q][6];
    mem_in_0[8*bw-1:7*bw] = K[q][7];
    mem_in_0[9*bw-1:8*bw] = K[q][8];
    mem_in_0[10*bw-1:9*bw] = K[q][9];
    mem_in_0[11*bw-1:10*bw] = K[q][10];
    mem_in_0[12*bw-1:11*bw] = K[q][11];
    mem_in_0[13*bw-1:12*bw] = K[q][12];
    mem_in_0[14*bw-1:13*bw] = K[q][13];
    mem_in_0[15*bw-1:14*bw] = K[q][14];
    mem_in_0[16*bw-1:15*bw] = K[q][15];

    #0.5 clk = 1'b1;  

  end

  #0.5 clk = 1'b0;  
  kmem_wr = 0;  
  qkmem_add = 0;
  #0.5 clk = 1'b1;  

  for (q=0; q<2; q=q+1) begin
    #0.5 clk = 1'b0;  
    #0.5 clk = 1'b1;   
  end


  for (q=col/2; q<col; q=q+1) begin

    #0.5 clk = 1'b0;  
    kmem_wr = 1; if (q>8) qkmem_add = qkmem_add + 1; 
    
    mem_in_1[1*bw-1:0*bw] = K[q][0];
    mem_in_1[2*bw-1:1*bw] = K[q][1];
    mem_in_1[3*bw-1:2*bw] = K[q][2];
    mem_in_1[4*bw-1:3*bw] = K[q][3];
    mem_in_1[5*bw-1:4*bw] = K[q][4];
    mem_in_1[6*bw-1:5*bw] = K[q][5];
    mem_in_1[7*bw-1:6*bw] = K[q][6];
    mem_in_1[8*bw-1:7*bw] = K[q][7];
    mem_in_1[9*bw-1:8*bw] = K[q][8];
    mem_in_1[10*bw-1:9*bw] = K[q][9];
    mem_in_1[11*bw-1:10*bw] = K[q][10];
    mem_in_1[12*bw-1:11*bw] = K[q][11];
    mem_in_1[13*bw-1:12*bw] = K[q][12];
    mem_in_1[14*bw-1:13*bw] = K[q][13];
    mem_in_1[15*bw-1:14*bw] = K[q][14];
    mem_in_1[16*bw-1:15*bw] = K[q][15];

    #0.5 clk = 1'b1;  

  end


  #0.5 clk = 1'b0;  
  kmem_wr = 0;  
  qkmem_add = 0;
  #0.5 clk = 1'b1;  
///////////////////////////////////////////



  for (q=0; q<2; q=q+1) begin
    #0.5 clk = 1'b0;  
    #0.5 clk = 1'b1;   
  end




/////  K data loading  /////
$display("##### K data loading to processor #####");

  for (q=0; q<(col/2)+1; q=q+1) begin
    #0.5 clk = 1'b0;  
    load = 1; 
    if (q==1) kmem_rd = 1;
    if (q>1) begin
       qkmem_add = qkmem_add + 1;
    end

    #0.5 clk = 1'b1;  
  end

  #0.5 clk = 1'b0;  
  kmem_rd = 0; qkmem_add = 0;
  #0.5 clk = 1'b1;  

  #0.5 clk = 1'b0;  
  load = 0; 
  #0.5 clk = 1'b1;  

///////////////////////////////////////////

 for (q=0; q<10; q=q+1) begin
    #0.5 clk = 1'b0;   
    #0.5 clk = 1'b1;   
 end





///// execution  /////
$display("##### execute #####");

  for (q=0; q<total_cycle; q=q+1) begin
    #0.5 clk = 1'b0;  
    execute = 1; 
    qmem_rd = 1;

    if (q>0) begin
       qkmem_add = qkmem_add + 1;
    end

    #0.5 clk = 1'b1;  
  end

  #0.5 clk = 1'b0;  
  qmem_rd = 0; qkmem_add = 0; execute = 0;
  #0.5 clk = 1'b1;  


///////////////////////////////////////////

 for (q=0; q<10; q=q+1) begin
    #0.5 clk = 1'b0;   
    #0.5 clk = 1'b1;   
 end

////////////// output fifo rd and wb to psum mem ///////////////////

$display("##### move ofifo to pmem #####");

  for (q=0; q<total_cycle; q=q+1) begin
    #0.5 clk = 1'b0;  
    ofifo_rd = 1; 
    pmem_wr = 1; 

    if (q>0) begin
       pmem_add = pmem_add + 1;
    end

    #0.5 clk = 1'b1;  
  end

  #0.5 clk = 1'b0;  
  pmem_wr = 0; pmem_add = 0; ofifo_rd = 0;
  #0.5 clk = 1'b1;  

///////////////////////////////////////////

 for (q=0; q<10; q=q+1) begin
    #0.5 clk = 1'b0;   
    #0.5 clk = 1'b1;   
 end

////////////////// move from pmem to sfp and process ////////////////////
  $display("#########Starting movement from pmem to sfp and processing#########");
  
  for(q=0;q<total_cycle*2;q=q+1) begin
    #0.5 clk = 1'b0;
    pmem_rd = 1;
    // ofifo_rd  =1;
    
    if(q%2==1) begin
        acc0 = 1;
        acc1 = 1;
    end
    else begin
	    acc0 = 0;
      acc1 = 0;
    end

    if(q>0 && q%2==0) begin
      pmem_add = pmem_add + 1;
    end
    #0.5 clk = 1'b1;


  end

  #0.5 clk = 1'b0;  
  pmem_rd = 0; ofifo_rd = 0; pmem_add = 0; acc0 = 0; acc1 = 0;
 
  #0.5 clk = 1'b1;


  #0.5 clk = 1'b0;
  #0.5 clk = 1'b1;
  #0.5 clk = 1'b0;
  #0.5 clk = 1'b1;


  for (q=0; q<total_cycle * 9; q=q+1) begin
    #0.5 clk = 1'b0;
    if(q%9 == 0) begin
      pmem_rd = 1;
    end
    
    if(q%9 == 1) begin
      canRead_0 = 1;
      canRead_1 = 1;
    end

    if(q%9 == 2) begin
      canRead_0 = 0;
      canRead_1 = 0;
    end

    if (q%9 == 6)begin
    div0 = 1;
    div1 = 1;
    end
    else begin
      div0 = 0;
      div1 = 0;
    end

   if (q%9 == 8)
    pmem_wr = 1;
   else
    pmem_wr = 0;


   if (q>0 && q%9 == 0) begin
    pmem_add = pmem_add + 1;
   end

    #0.5 clk = 1'b1;
  end

  #0.5 clk = 1'b0;  
  pmem_rd = 0; pmem_add = 0; div0 = 0; div1 = 0;
  #0.5 clk = 1'b1;

  // for(q=0;q<total_cycle+2;q=q+1) begin
  //   #0.5 clk = 1'b0;
  //   fifo_ext_rd = 1'b1;
    
  //   fifo_out[q] = sum_out;
  //   #0.5 clk = 1'b1;
  // end

  #10 $finish;


end

endmodule



